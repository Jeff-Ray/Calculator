/********************************************************************
*                      二进制转BCD（左移加三算法）
*    说明： 如果某一权位（百位，十位，个位）大于或者等于5，那么此权位加3。
*          将二进制数，左移1位到BCD移位寄存器中。
*          如果二进制数据位都移动完毕，计算结束
*	功能：将二进制码转为十进制BCD码
*	作者：Ray
*	起始时间：2021-4-24
*	完成时间：2021-5-26
********************************************************************/
module bcd_d(

		input wire [13:0] binary,
		output wire [3:0] g,
		output wire [3:0] s,
		output wire [3:0] b,
		output wire [3:0] q
	
    	);

    reg [29:0] z;

    always @ (*)
    begin
        z = 29'b0;                           //置 0
        z[13:0] = binary;                     //读入低 8 位
        repeat (14)                            //重复 8 次
        begin
            if(z[17:14]>4)                   //大于 4 就加 3
               z[17:14] = z[17:14] + 2'b11;
            if(z[21:18]>4)
               z[21:18] = z[21:18] + 2'b11;
				if(z[25:22]>4)
               z[25:22] = z[25:22] + 2'b11;
				if(z[29:26]>4)
               z[29:26] = z[29:26] + 2'b11;
            z[29:1] = z[28:0];               //左移一位
			end
		end

        //输出 BCD码
        assign q = z[29:26]; 
		assign b = z[25:22];                     
		assign s = z[21:18];
		assign g = z[17:14];
    
endmodule
